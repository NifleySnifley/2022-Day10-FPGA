
module ROM (
	input wire [addr_bits-1:0] addr,
	output reg [data_width-1:0] data,  // reg (not wire)
	output wire [7:0] screen_w,
	output wire [7:0] screen_h
);
parameter addr_bits = 8,
		  data_width = 8;

assign screen_w = 8'd40;
assign screen_h = 8'd6;

always_comb
begin
	case(addr)
		8'd0 : data = 0;
		8'd1 : data = 2;
		8'd2 : data = 0;
		8'd3 : data = 3;
		8'd4 : data = 0;
		8'd5 : data = 0;
		8'd6 : data = 0;
		8'd7 : data = 1;
		8'd8 : data = 0;
		8'd9 : data = 5;
		8'd10 : data = 0;
		8'd11 : data = -1;
		8'd12 : data = 0;
		8'd13 : data = 5;
		8'd14 : data = 0;
		8'd15 : data = 1;
		8'd16 : data = 0;
		8'd17 : data = 0;
		8'd18 : data = 0;
		8'd19 : data = 4;
		8'd20 : data = 0;
		8'd21 : data = 0;
		8'd22 : data = 0;
		8'd23 : data = 5;
		8'd24 : data = 0;
		8'd25 : data = -5;
		8'd26 : data = 0;
		8'd27 : data = 6;
		8'd28 : data = 0;
		8'd29 : data = 3;
		8'd30 : data = 0;
		8'd31 : data = 1;
		8'd32 : data = 0;
		8'd33 : data = 5;
		8'd34 : data = 0;
		8'd35 : data = 1;
		8'd36 : data = 0;
		8'd37 : data = 0;
		8'd38 : data = -38;
		8'd39 : data = 0;
		8'd40 : data = 41;
		8'd41 : data = 0;
		8'd42 : data = -22;
		8'd43 : data = 0;
		8'd44 : data = -14;
		8'd45 : data = 0;
		8'd46 : data = 7;
		8'd47 : data = 0;
		8'd48 : data = 0;
		8'd49 : data = 0;
		8'd50 : data = 3;
		8'd51 : data = 0;
		8'd52 : data = -2;
		8'd53 : data = 0;
		8'd54 : data = 2;
		8'd55 : data = 0;
		8'd56 : data = 0;
		8'd57 : data = 17;
		8'd58 : data = 0;
		8'd59 : data = -12;
		8'd60 : data = 0;
		8'd61 : data = 5;
		8'd62 : data = 0;
		8'd63 : data = 2;
		8'd64 : data = 0;
		8'd65 : data = -16;
		8'd66 : data = 0;
		8'd67 : data = 17;
		8'd68 : data = 0;
		8'd69 : data = 2;
		8'd70 : data = 0;
		8'd71 : data = 5;
		8'd72 : data = 0;
		8'd73 : data = 2;
		8'd74 : data = 0;
		8'd75 : data = -30;
		8'd76 : data = 0;
		8'd77 : data = 0;
		8'd78 : data = -6;
		8'd79 : data = 0;
		8'd80 : data = 1;
		8'd81 : data = 0;
		8'd82 : data = 0;
		8'd83 : data = 5;
		8'd84 : data = 0;
		8'd85 : data = 0;
		8'd86 : data = 0;
		8'd87 : data = 0;
		8'd88 : data = 5;
		8'd89 : data = 0;
		8'd90 : data = -12;
		8'd91 : data = 0;
		8'd92 : data = 17;
		8'd93 : data = 0;
		8'd94 : data = 0;
		8'd95 : data = 0;
		8'd96 : data = 0;
		8'd97 : data = 0;
		8'd98 : data = 5;
		8'd99 : data = 0;
		8'd100 : data = 10;
		8'd101 : data = 0;
		8'd102 : data = -9;
		8'd103 : data = 0;
		8'd104 : data = 2;
		8'd105 : data = 0;
		8'd106 : data = 5;
		8'd107 : data = 0;
		8'd108 : data = 2;
		8'd109 : data = 0;
		8'd110 : data = -5;
		8'd111 : data = 0;
		8'd112 : data = 6;
		8'd113 : data = 0;
		8'd114 : data = 4;
		8'd115 : data = 0;
		8'd116 : data = 0;
		8'd117 : data = 0;
		8'd118 : data = -37;
		8'd119 : data = 0;
		8'd120 : data = 0;
		8'd121 : data = 0;
		8'd122 : data = 17;
		8'd123 : data = 0;
		8'd124 : data = -12;
		8'd125 : data = 0;
		8'd126 : data = 30;
		8'd127 : data = 0;
		8'd128 : data = -23;
		8'd129 : data = 0;
		8'd130 : data = 2;
		8'd131 : data = 0;
		8'd132 : data = 0;
		8'd133 : data = 3;
		8'd134 : data = 0;
		8'd135 : data = -17;
		8'd136 : data = 0;
		8'd137 : data = 22;
		8'd138 : data = 0;
		8'd139 : data = 0;
		8'd140 : data = 0;
		8'd141 : data = 0;
		8'd142 : data = 5;
		8'd143 : data = 0;
		8'd144 : data = 0;
		8'd145 : data = -10;
		8'd146 : data = 0;
		8'd147 : data = 11;
		8'd148 : data = 0;
		8'd149 : data = 4;
		8'd150 : data = 0;
		8'd151 : data = 0;
		8'd152 : data = 5;
		8'd153 : data = 0;
		8'd154 : data = -2;
		8'd155 : data = 0;
		8'd156 : data = 0;
		8'd157 : data = -6;
		8'd158 : data = 0;
		8'd159 : data = -29;
		8'd160 : data = 0;
		8'd161 : data = 37;
		8'd162 : data = 0;
		8'd163 : data = -30;
		8'd164 : data = 0;
		8'd165 : data = 27;
		8'd166 : data = 0;
		8'd167 : data = -2;
		8'd168 : data = 0;
		8'd169 : data = -22;
		8'd170 : data = 0;
		8'd171 : data = 0;
		8'd172 : data = 3;
		8'd173 : data = 0;
		8'd174 : data = 2;
		8'd175 : data = 0;
		8'd176 : data = 0;
		8'd177 : data = 7;
		8'd178 : data = 0;
		8'd179 : data = -2;
		8'd180 : data = 0;
		8'd181 : data = 2;
		8'd182 : data = 0;
		8'd183 : data = 5;
		8'd184 : data = 0;
		8'd185 : data = -5;
		8'd186 : data = 0;
		8'd187 : data = 6;
		8'd188 : data = 0;
		8'd189 : data = 2;
		8'd190 : data = 0;
		8'd191 : data = 2;
		8'd192 : data = 0;
		8'd193 : data = 5;
		8'd194 : data = 0;
		8'd195 : data = -25;
		8'd196 : data = 0;
		8'd197 : data = 0;
		8'd198 : data = -10;
		8'd199 : data = 0;
		8'd200 : data = 0;
		8'd201 : data = 1;
		8'd202 : data = 0;
		8'd203 : data = 0;
		8'd204 : data = 2;
		8'd205 : data = 0;
		8'd206 : data = 0;
		8'd207 : data = 0;
		8'd208 : data = 0;
		8'd209 : data = 0;
		8'd210 : data = 7;
		8'd211 : data = 0;
		8'd212 : data = 1;
		8'd213 : data = 0;
		8'd214 : data = 4;
		8'd215 : data = 0;
		8'd216 : data = 1;
		8'd217 : data = 0;
		8'd218 : data = 0;
		8'd219 : data = 2;
		8'd220 : data = 0;
		8'd221 : data = 0;
		8'd222 : data = 3;
		8'd223 : data = 0;
		8'd224 : data = 5;
		8'd225 : data = 0;
		8'd226 : data = -1;
		8'd227 : data = 0;
		8'd228 : data = 0;
		8'd229 : data = 3;
		8'd230 : data = 0;
		8'd231 : data = 5;
		8'd232 : data = 0;
		8'd233 : data = 2;
		8'd234 : data = 0;
		8'd235 : data = 1;
		8'd236 : data = 0;
		8'd237 : data = 0;
		8'd238 : data = 0;
		8'd239 : data = 0;
		default : data = 8'b00000000;
	endcase 
end

endmodule
